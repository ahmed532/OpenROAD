module SoC (
    input clk,
    input rst,
    inout [31:0] data_bus
);
endmodule
