module TopDesign (
  input clk,
  input reset
);
endmodule
